
module clock_manual (
    input button,
	 output clk
);

	assign clk = button;
 
    
endmodule

